library ieee;
use IEEE.std_Logic_1164.all;
use IEEE.NUMERIC_STD.ALL; 
use IEEE.std_Logic_unsigned.all;
use work.V1495_regs.all;
use work.functions.all;
entity V1495_regs_communication is
  generic(
    N_R_REGS : integer := 18;
    N_RW_REGS : integer := 84
  );
  port(
    -- Data clock
    clk_data   : in std_logic;
    -- Local Bus in/out signals
    nLBRES     : in     std_logic;
    nBLAST     : in     std_logic;
    WnR        : in     std_logic;
    nADS       : in     std_logic;
    LCLK       : in     std_logic;
    nREADY     : out    std_logic;
    nINT       : out    std_logic;
    LAD        : inout  std_logic_vector(15 DOWNTO 0);
    ADDR_W : out std_logic_vector(11 downto 0);
    REG_R  : in reg_data(N_R_REGS - 1 downto 0);
    REG_RW : out reg_data(N_RW_REGS - 1 downto 0)
  );
end V1495_regs_communication;
architecture rtl of V1495_regs_communication is
begin
  ADDR_W <= x"000";
  REG_RW(0) <= x"00000000";
  REG_RW(1) <= x"00000000";
  REG_RW(2) <= x"00000000";
  REG_RW(3) <= x"00000000";
  REG_RW(4) <= x"00000000";
  REG_RW(5) <= x"00000000";
  REG_RW(6) <= x"0a0a0a0a";
  REG_RW(7) <= x"0a0a0a08";
  REG_RW(8) <= x"00000000";
  REG_RW(9) <= x"00000000";
  REG_RW(10) <= x"00000000";
  REG_RW(11) <= x"00000000";
  REG_RW(12) <= x"00000000";
  REG_RW(13) <= x"00000000";
  REG_RW(14) <= x"00000000";
  REG_RW(15) <= x"00000000";
  REG_RW(16) <= x"00000000";
  REG_RW(17) <= x"00000000";
  REG_RW(18) <= x"00000000";
  REG_RW(19) <= x"00000000";
  REG_RW(20) <= x"00000000";
  REG_RW(21) <= x"00000000";
  REG_RW(22) <= x"05050505";
  REG_RW(23) <= x"05050505";
  REG_RW(24) <= x"00000000";
  REG_RW(25) <= x"00000000";
  REG_RW(26) <= x"00000000";
  REG_RW(27) <= x"00000000";
  REG_RW(28) <= x"00000000";
  REG_RW(29) <= x"00000000";
  REG_RW(30) <= x"00000000";
  REG_RW(31) <= x"00000000";
  REG_RW(32) <= x"00000000";
  REG_RW(33) <= x"00000000";
  REG_RW(34) <= x"00000000";
  REG_RW(35) <= x"00000000";
  REG_RW(36) <= x"00000000";
  REG_RW(37) <= x"00000000";
  REG_RW(38) <= x"00000000";
  REG_RW(39) <= x"00000000";
  REG_RW(40) <= x"00000000";
  REG_RW(41) <= x"00000000";
  REG_RW(42) <= x"00000000";
  REG_RW(43) <= x"00000000";
  REG_RW(44) <= x"00000000";
  REG_RW(45) <= x"00000000";
  REG_RW(46) <= x"00000000";
  REG_RW(47) <= x"00000000";
  REG_RW(48) <= x"00000000";
  REG_RW(49) <= x"00000000";
  REG_RW(50) <= x"00000000";
  REG_RW(51) <= x"00000000";
  REG_RW(52) <= x"00000000";
  REG_RW(53) <= x"00000000";
  REG_RW(54) <= x"00000050";
  REG_RW(55) <= x"00000000";
  REG_RW(56) <= x"00000000";
  REG_RW(57) <= x"00000000";
  REG_RW(58) <= x"00000000";
  REG_RW(59) <= x"00000000";
  REG_RW(60) <= x"00000000";
  REG_RW(61) <= x"00000000";
  REG_RW(62) <= x"00000000";
  REG_RW(63) <= x"00000000";
  REG_RW(64) <= x"00000000";
  REG_RW(65) <= x"00000000";
  REG_RW(66) <= x"00000000";
  REG_RW(67) <= x"00000000";
  REG_RW(68) <= x"00000000";
  REG_RW(69) <= x"00000000";
  REG_RW(70) <= x"00000000";
  REG_RW(71) <= x"00000000";
  REG_RW(72) <= x"00000000";
  REG_RW(73) <= x"00000000";
  REG_RW(74) <= x"0000000e";
  REG_RW(75) <= x"00000000";
  REG_RW(76) <= x"00000000";
  REG_RW(77) <= x"0000000f";
  REG_RW(78) <= x"00000000";
  REG_RW(79) <= x"00000000";
  REG_RW(80) <= x"00000000";
  REG_RW(81) <= x"00000000";
  REG_RW(82) <= x"00000000";
  REG_RW(83) <= x"00000000";
  REG_RW(84) <= x"00000000";
  REG_RW(85) <= x"00000000";
  REG_RW(86) <= x"00000000";
  REG_RW(87) <= x"00000000";
  REG_RW(88) <= x"00000000";
  REG_RW(89) <= x"00000001";
  REG_RW(90) <= x"00000000";
  REG_RW(91) <= x"00000000";
  REG_RW(92) <= x"00000060";
  REG_RW(93) <= x"000000e0";
  REG_RW(94) <= x"0000006b";
  REG_RW(95) <= x"000000ec";
  REG_RW(96) <= x"00000084";
  REG_RW(97) <= x"00000085";
  REG_RW(98) <= x"00000086";
  REG_RW(99) <= x"00000087";
  REG_RW(100) <= x"00000000";
  REG_RW(101) <= x"00000000";
  REG_RW(102) <= x"00000000";
  REG_RW(103) <= x"00000000";
  REG_RW(104) <= x"00000000";
  REG_RW(105) <= x"00000000";
  REG_RW(106) <= x"00000000";
  REG_RW(107) <= x"00000000";
  REG_RW(108) <= x"00000000";
  REG_RW(109) <= x"00000000";
  REG_RW(110) <= x"00000000";
  REG_RW(111) <= x"00003332";
  REG_RW(112) <= x"00000000";
  REG_RW(113) <= x"00000000";
  REG_RW(114) <= x"00000000";
  REG_RW(115) <= x"00000000";
  REG_RW(116) <= x"00000000";
  REG_RW(117) <= x"00000000";
  REG_RW(118) <= x"00000000";
  REG_RW(119) <= x"00000000";
  REG_RW(120) <= x"00000000";
  REG_RW(121) <= x"00000000";
  REG_RW(122) <= x"00000000";
  REG_RW(123) <= x"00000000";
  REG_RW(124) <= x"00000000";
  REG_RW(125) <= x"00000000";
  REG_RW(126) <= x"00000000";
  REG_RW(127) <= x"00000000";
  REG_RW(128) <= x"00000000";
  REG_RW(129) <= x"00000000";
  REG_RW(130) <= x"00000000";
  REG_RW(131) <= x"00000000";
  REG_RW(132) <= x"00000000";
  REG_RW(133) <= x"00000000";
  REG_RW(134) <= x"00000001";
  REG_RW(135) <= x"00000000";
  REG_RW(136) <= x"00000000";
  REG_RW(137) <= x"00000000";
  REG_RW(138) <= x"00000000";
  REG_RW(139) <= x"00000000";
  REG_RW(140) <= x"00000000";
  REG_RW(141) <= x"00000000";
  REG_RW(142) <= x"00000000";
  REG_RW(143) <= x"00000000";
  REG_RW(144) <= x"00000010";
  REG_RW(145) <= x"00000000";
  REG_RW(146) <= x"00000000";
  REG_RW(147) <= x"00000000";
  REG_RW(148) <= x"00000000";
  REG_RW(149) <= x"00000000";
  REG_RW(150) <= x"00000000";
  REG_RW(151) <= x"00000000";
  REG_RW(152) <= x"00000000";
  REG_RW(153) <= x"00000000";
  REG_RW(154) <= x"00000000";
end architecture rtl;
